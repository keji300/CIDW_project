`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/01/12 17:22:51
// Design Name: 
// Module Name: decode7_80
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module decode7_80(
input [6:0] a,
output reg [79:0]b
    );
    always @ (*)
    begin
    	case (a)
    	0  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001;
    	1  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010;
    	2  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100;
    	3  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000;
    	4  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000;
    	5  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000;
    	6  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000;
    	7  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000;
    	8  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000;
    	9  : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000;
    	10 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000;
    	11 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000;
    	12 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000;
    	13 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
    	14 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000;
    	15 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000;
    	16 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000;
    	17 : b <= 80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000;
    	18 : b <= 80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000;
    	19 : b <= 80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000;
    	20 : b <= 80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000;
    	21 : b <= 80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000;
    	22 : b <= 80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000;
    	23 : b <= 80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000;
    	24 : b <= 80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000;
    	25 : b <= 80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000;
    	26 : b <= 80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000;
    	27 : b <= 80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000;
    	28 : b <= 80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000;
    	29 : b <= 80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000;
    	30 : b <= 80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000;
    	31 : b <= 80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000;
    	32 : b <= 80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000;
    	33 : b <= 80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000;
    	34 : b <= 80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000;
    	35 : b <= 80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000;
    	36 : b <= 80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000;
    	37 : b <= 80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000;
    	38 : b <= 80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000;
    	39 : b <= 80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000;
    	40 : b <= 80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000;
    	41 : b <= 80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000;
    	42 : b <= 80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000;
    	43 : b <= 80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000;
    	44 : b <= 80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000;
    	45 : b <= 80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000;
    	46 : b <= 80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000;
    	47 : b <= 80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000;
    	48 : b <= 80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000;
    	49 : b <= 80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000;
    	50 : b <= 80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000;
    	51 : b <= 80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000;
    	52 : b <= 80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000;
    	53 : b <= 80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000;
    	54 : b <= 80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000;
    	55 : b <= 80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000;
    	56 : b <= 80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000;
    	57 : b <= 80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000;
    	58 : b <= 80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000;
    	59 : b <= 80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000;
    	60 : b <= 80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000;
    	61 : b <= 80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000;
    	62 : b <= 80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000;
    	63 : b <= 80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000;
    	64 : b <= 80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000;
    	65 : b <= 80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000;
    	66 : b <= 80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000;
    	67 : b <= 80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000;
    	68 : b <= 80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000;
    	69 : b <= 80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000;
    	70 : b <= 80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000;
    	71 : b <= 80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000;
    	72 : b <= 80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000;
    	73 : b <= 80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000;
    	74 : b <= 80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000;
    	75 : b <= 80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000;
    	76 : b <= 80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000;
    	77 : b <= 80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000;
    	78 : b <= 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000;
    	79 : b <= 80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000;
		default: b <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    	endcase
    end
    
    
    
    
endmodule
